module DoubleDabble();
endmodule