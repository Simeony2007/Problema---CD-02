modulo main();


	Multiplicador mult1(S, A, B, Clock)


endmodule