module RPNInput(S, A, FF0, FF1, FF2, FF3, Contador);
	input A, FF0, FF1, FF2, FF3;
	input [1:0]Contador;
	output [3:0]S;
	wire [3:0]T;

	
	
endmodule