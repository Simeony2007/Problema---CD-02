module Multiplicador();

	// Trabalhando

endmodule