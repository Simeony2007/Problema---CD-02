//============================================================
// BINÁRIO (8 bits) -> 3 DISPLAYS OCTAL ============================================================
module ConversorOctal(
    input  [7:0] BIN,
    output [2:0] A, B, C, D, E, F, G
);

    // -------------------------
    // DIGITO menos significativo (O0)
    // -------------------------
    wire [2:0] O0 = BIN[2:0];

    // -------------------------
    // DIGITO do meio (O1)
    // -------------------------
    wire [2:0] O1 = BIN[5:3];

    // -------------------------
    // DIGITO mais significativo (O2) - totalmente estrutural
    // -------------------------
    wire O2_2, O2_1, O2_0;
    // Bits altos da entrada
    and (O2_2, BIN[7], 1'b1); // simplesmente BIN[7]
    and (O2_1, BIN[6], 1'b1); // simplesmente BIN[6]
    wire zero;
    and (O2_0, 1'b0, 1'b0);   // bit menos significativo sempre 0 (GND)

    // -------------------------
    // DIGITO 0 (O0)
    // -------------------------
    not (n0_2, O0[2]);
    not (n0_1, O0[1]);
    not (n0_0, O0[0]);

    wire m0_0, m0_1, m0_2, m0_3, m0_4, m0_5, m0_6, m0_7;
    and (m0_0, n0_2, n0_1, n0_0);
    and (m0_1, n0_2, n0_1, O0[0]);
    and (m0_2, n0_2, O0[1], n0_0);
    and (m0_3, n0_2, O0[1], O0[0]);
    and (m0_4, O0[2], n0_1, n0_0);
    and (m0_5, O0[2], n0_1, O0[0]);
    and (m0_6, O0[2], O0[1], n0_0);
    and (m0_7, O0[2], O0[1], O0[0]);

    or (A[0], m0_0,m0_2,m0_3,m0_5,m0_6,m0_7);
    or (B[0], m0_1,m0_2,m0_3,m0_4,m0_7);
    or (C[0], m0_1,m0_3,m0_5,m0_6,m0_7);
    or (D[0], m0_0,m0_2,m0_3,m0_5,m0_6,m0_7);
    or (E[0], m0_0,m0_2,m0_6);
    or (F[0], m0_0,m0_4,m0_5,m0_6,m0_7);
    or (G[0], m0_2,m0_3,m0_4,m0_5,m0_6,m0_7);

    // -------------------------
    // DIGITO 1 (O1)
    // -------------------------
    not (n1_2, O1[2]);
    not (n1_1, O1[1]);
    not (n1_0, O1[0]);

    wire m1_0, m1_1, m1_2, m1_3, m1_4, m1_5, m1_6, m1_7;
    and (m1_0, n1_2,n1_1,n1_0);
    and (m1_1, n1_2,n1_1,O1[0]);
    and (m1_2, n1_2,O1[1],n1_0);
    and (m1_3, n1_2,O1[1],O1[0]);
    and (m1_4, O1[2],n1_1,n1_0);
    and (m1_5, O1[2],n1_1,O1[0]);
    and (m1_6, O1[2],O1[1],n1_0);
    and (m1_7, O1[2],O1[1],O1[0]);

    or (A[1], m1_0,m1_2,m1_3,m1_5,m1_6,m1_7);
    or (B[1], m1_1,m1_2,m1_3,m1_4,m1_7);
    or (C[1], m1_1,m1_3,m1_5,m1_6,m1_7);
    or (D[1], m1_0,m1_2,m1_3,m1_5,m1_6,m1_7);
    or (E[1], m1_0,m1_2,m1_6);
    or (F[1], m1_0,m1_4,m1_5,m1_6,m1_7);
    or (G[1], m1_2,m1_3,m1_4,m1_5,m1_6,m1_7);

    // -------------------------
    // DIGITO 2 (O2)
    // -------------------------
    not (n2_2, O2_2);
    not (n2_1, O2_1);
    not (n2_0, O2_0);

    wire m2_0, m2_1, m2_2, m2_3, m2_4, m2_5, m2_6, m2_7;
    and (m2_0, n2_2,n2_1,n2_0);
    and (m2_1, n2_2,n2_1,O2_0);
    and (m2_2, n2_2,O2_1,n2_0);
    and (m2_3, n2_2,O2_1,O2_0);
    and (m2_4, O2_2,n2_1,n2_0);
    and (m2_5, O2_2,n2_1,O2_0);
    and (m2_6, O2_2,O2_1,n2_0);
    and (m2_7, O2_2,O2_1,O2_0);

    or (A[2], m2_0,m2_2,m2_3,m2_5,m2_6,m2_7);
    or (B[2], m2_1,m2_2,m2_3,m2_4,m2_7);
    or (C[2], m2_1,m2_3,m2_5,m2_6,m2_7);
    or (D[2], m2_0,m2_2,m2_3,m2_5,m2_6,m2_7);
    or (E[2], m2_0,m2_2,m2_6);
    or (F[2], m2_0,m2_4,m2_5,m2_6,m2_7);
    or (G[2], m2_2,m2_3,m2_4,m2_5,m2_6,m2_7);

endmodule
