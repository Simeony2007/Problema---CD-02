module SomComp8bits(S, Cout, A, B, Cin);
	// DECLARANDO ENTRADAS, SAIDAS E FIOS:
	input [7:0]A;
	input [7:0]B;
	input Cin;
	output [7:0]S;
	output Cout;
	wire [6:0]T;
	
	// INSTANCIAÇÃO DO SOMADOR COMPLETO DE 1 BIT:
	SomComp1bit U0(S[0], T[0], A[0], B[0], Cin);
	SomComp1bit U1(S[1], T[1], A[1], B[1], T[0]);
	SomComp1bit U2(S[2], T[2], A[2], B[2], T[1]);
	SomComp1bit U3(S[3], T[3], A[3], B[3], T[2]);
	SomComp1bit U4(S[4], T[4], A[4], B[4], T[3]);
	SomComp1bit U5(S[5], T[5], A[5], B[5], T[4]);
	SomComp1bit U6(S[6], T[6], A[6], B[6], T[5]);
	SomComp1bit U7(S[7], Cout, A[7], B[7], T[6]);
	
endmodule