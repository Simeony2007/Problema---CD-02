module Multiplicador(S, A, B, Clock, Cont);
	input [7:0]A;
	input [7:0]B;
	input Clock;
	input Cont;
	output [15:0]S;
	wire [7:0]R;
	wire [7:0]T;
	
	
	

endmodule