module FlipFlop(Out, Set, Reset);

	reg

endmodule