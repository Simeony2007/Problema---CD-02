module MUX_16bit_8para1(Y, S, I0, I1, I2, I3, I4, I5, I6, I7);
    output [15:0] Y;
    input  [2:0] S;
    input  [15:0] I0, I1, I2, I3, I4, I5, I6, I7;

    // Instancia 16 MUXes de 1 bit
    MUX_1bit_8para1 m0(Y[0], {I7[0],I6[0],I5[0],I4[0],I3[0],I2[0],I1[0],I0[0]}, S);
    MUX_1bit_8para1 m1(Y[1], {I7[1],I6[1],I5[1],I4[1],I3[1],I2[1],I1[1],I0[1]}, S);
    MUX_1bit_8para1 m2(Y[2], {I7[2],I6[2],I5[2],I4[2],I3[2],I2[2],I1[2],I0[2]}, S);
    MUX_1bit_8para1 m3(Y[3], {I7[3],I6[3],I5[3],I4[3],I3[3],I2[3],I1[3],I0[3]}, S);
    MUX_1bit_8para1 m4(Y[4], {I7[4],I6[4],I5[4],I4[4],I3[4],I2[4],I1[4],I0[4]}, S);
    MUX_1bit_8para1 m5(Y[5], {I7[5],I6[5],I5[5],I4[5],I3[5],I2[5],I1[5],I0[5]}, S);
    MUX_1bit_8para1 m6(Y[6], {I7[6],I6[6],I5[6],I4[6],I3[6],I2[6],I1[6],I0[6]}, S);
    MUX_1bit_8para1 m7(Y[7], {I7[7],I6[7],I5[7],I4[7],I3[7],I2[7],I1[7],I0[7]}, S);
    MUX_1bit_8para1 m8(Y[8], {I7[8],I6[8],I5[8],I4[8],I3[8],I2[8],I1[8],I0[8]}, S);
    MUX_1bit_8para1 m9(Y[9], {I7[9],I6[9],I5[9],I4[9],I3[9],I2[9],I1[9],I0[9]}, S);
    MUX_1bit_8para1 m10(Y[10], {I7[10],I6[10],I5[10],I4[10],I3[10],I2[10],I1[10],I0[10]}, S);
    MUX_1bit_8para1 m11(Y[11], {I7[11],I6[11],I5[11],I4[11],I3[11],I2[11],I1[11],I0[11]}, S);
    MUX_1bit_8para1 m12(Y[12], {I7[12],I6[12],I5[12],I4[12],I3[12],I2[12],I1[12],I0[12]}, S);
    MUX_1bit_8para1 m13(Y[13], {I7[13],I6[13],I5[13],I4[13],I3[13],I2[13],I1[13],I0[13]}, S);
    MUX_1bit_8para1 m14(Y[14], {I7[14],I6[14],I5[14],I4[14],I3[14],I2[14],I1[14],I0[14]}, S);
    MUX_1bit_8para1 m15(Y[15], {I7[15],I6[15],I5[15],I4[15],I3[15],I2[15],I1[15],I0[15]}, S);
endmodule